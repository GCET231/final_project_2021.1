////////////////////////////////////////
// Projeto Final 2021.1
// João Bittencourt
////////////////////////////////////////
// Como tenho um coração muito grande e magnânimo, deixo aqui uma parte do módulo do Black Jack (\o/)

module BlackJackFSM (
   input CLK, 
   input RESET, 
   input STAY, 
   input HIT, 
   input [3:0] CARD, 
   output WIN, 
   output LOSE, 
   output TIE, 
   // Sinais para controle de envio de cartas para o Dealer
   // usados apenas para depuração no test bench.
   output DHIT,  
   output DSTAY
);

// FSM States

// Internal Signals

// Current State

// Next State Logic

// Output Logic

endmodule